/*Array Manipulation methods:it provides several built in methods to operate on arrays
1.Array ordering methods
2.Array reduction methods
3.Array locator method
4.Array iterator index querying


1.Array ordering methods:
it operates on 1d arrays or queues
these methods useful for reordering the array elements
built in array ordering methods are:
a)reverse
b)sort
c)rsort
d)shuffle*/
//we cant apply array ordering methods to associative arrays